library verilog;
use verilog.vl_types.all;
entity tb_ahb_lite is
end tb_ahb_lite;
