library verilog;
use verilog.vl_types.all;
entity tb_spi is
end tb_spi;
